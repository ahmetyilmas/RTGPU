`timescale 1ns/1ps

`include "Types.sv"
`include "Parameters.sv"


module RayCore #(
    parameter int WIDTH = 20,
    parameter int QBITS = 12
) (
    input clk,
    input reset,
    input start,
    input Cam_t camera_in
);

endmodule

`include "../Types.sv"
`include "../Parameters.sv"

module LambertianShader #(
    parameter int WIDTH = 20,
    parameter int Q_BITS = 12
)(
    input clk,
    input reset,
    input start,
    input Color_t color_in

);

endmodule
